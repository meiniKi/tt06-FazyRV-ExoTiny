(* blackbox *)
module sky130_fd_sc_hd__dlygate4sd3_1 (
  input   A,
  output  X
);

endmodule 